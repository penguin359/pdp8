localparam [2:0] OPCODE_AND = 3'b000;
localparam [2:0] OPCODE_TAD = 3'b001;
localparam [2:0] OPCODE_ISZ = 3'b010;
localparam [2:0] OPCODE_DCA = 3'b011;
localparam [2:0] OPCODE_JMS = 3'b100;
localparam [2:0] OPCODE_JMP = 3'b101;
localparam [2:0] OPCODE_IOT = 3'b110;
localparam [2:0] OPCODE_OPR = 3'b111;

localparam Z_BIT = 7;
localparam I_BIT = 8;

class uarttx_driver extends uvm_driver #(uarttx_transaction);
endclass: uarttx_driver
